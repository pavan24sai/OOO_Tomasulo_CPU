`ifndef MACROS_SVH
`define MACROS_SVH

`define BENCHMARK "test_add_sub" 	// test_add_sub | test_dependencies	| test_fibonacci | test_mem_simple | test_sb_simple | test_sb_type
`define SIM_CYCLES 685          	// change number of cycles to run simulation for
`define TESTING_NON_SYNTH       	// comment out to disable automated testing

`endif  // MACROS_SVH
